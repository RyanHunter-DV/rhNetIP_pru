module ncpc_arb (
); // {


endmodule // }
